module hazard(input  logic			MemtoRegE,
			  input  logic			RegWriteW,
			  input  logic			RegWriteM,
			  input  logic			Match,
			  output logic			ForwardAE,
			  output logic			ForwardBE,
			  output logic			FlushE,
			  output logic			StallD,
			  output logic			StallF);
	
	
	
endmodule
